`define DW 8
`define AW 8
