`include "apb_interface.sv"
`include "apb_sequence_item.sv"
`include "apb_sequence.sv"
`include "apb_sequencer.sv"
`include "apb_driver.sv"
`include "apb_in_mon.sv"
`include "apb_out_mon.sv"
`include "apb_active_agent.sv"
`include "apb_passive_agent.sv"
`include "apb_scoreboard.sv"
//`include "apb_coverage.sv"
`include "apb_env.sv"
`include "apb_test.sv"
